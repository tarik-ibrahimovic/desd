library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity balance_controller is
	generic (
		TDATA_WIDTH		: positive := 24;
		BALANCE_WIDTH	: positive := 10;
		BALANCE_STEP_2	: positive := 6		-- i.e., balance_values_per_step = 2**VOLUME_STEP_2
	);
	Port (
		aclk			: in std_logic;
		aresetn			: in std_logic;

		s_axis_tvalid	: in std_logic;
		s_axis_tdata	: in std_logic_vector(TDATA_WIDTH-1 downto 0);
		s_axis_tready	: out std_logic;
		s_axis_tlast	: in std_logic;

		m_axis_tvalid	: out std_logic;
		m_axis_tdata	: out std_logic_vector(TDATA_WIDTH-1 downto 0);
		m_axis_tready	: in std_logic;
		m_axis_tlast	: out std_logic;

		balance			: in std_logic_vector(BALANCE_WIDTH-1 downto 0)
	);
end balance_controller;

architecture Behavioral of balance_controller is
    signal N : natural range 0 to 2**BALANCE_WIDTH-1;   
    signal t_data : std_logic_vector(TDATA_WIDTH-1 downto 0);
    
begin
    
    N               <= to_integer(unsigned(balance(BALANCE_WIDTH-2 downto 0)) srl BALANCE_STEP_2); 
    t_data          <= s_axis_tdata when s_axis_tlast = balance(BALANCE_WIDTH-1) else std_logic_vector(signed(s_axis_tdata) srl N); 
    
end Behavioral;
